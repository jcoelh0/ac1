library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.DisplayUnit_pkg.all;

entity Ram is
	generic(	ADDR_BUS_SIZE 	: positive := 6;
				DATA_BUS_SIZE	: positive := 32);
	port(	clk 		: 	in 	std_logic;
			readEn	:	in		std_logic;
			writeEn	:	in		std_logic;
			address	:	in		std_logic_vector(ADDR_BUS_SIZE-1 downto 0);
			writeData:	in		std_logic_vector(DATA_BUS_SIZE-1 downto 0);
			readData	:	out	std_logic_vector(DATA_BUS_SIZE-1 downto 0));
end Ram;

architecture Behavioral of Ram is
	constant NUM_WORDS : positive := (2**ADDR_BUS_SIZE);
	subtype TData is std_logic_vector(DATA_BUS_SIZE-1 downto 0);
	type TMemory is array(0 to NUM_WORDS-1) of TData;
	signal s_memory : TMemory:= (	X"8c010000",	-- lw $1, 0x0000($0)
											X"20210004",	-- addi $1,$1,4
											X"AC010004",	-- sw $1, 4($0)
											others => X"00000000");

begin
	process(clk)
	begin
		if(rising_edge(clk)) then
			if(writeEn = '1') then
				s_memory(to_integer(unsigned(address))) <= writeData;
			end if;
		end if;
	end process;
	
	readData <= s_memory(to_integer(unsigned(address))) when
					(readEn = '1') else (others => '-');

	DU_DMdata <= s_memory(to_integer(unsigned(DU_DMaddr)));
end Behavioral;